//-----------------------------------------------------------------------------
// Title                 : random_tb
// Project               : ECE 411 mp_verif
//-----------------------------------------------------------------------------
// File                  : random_tb.sv
// Author                : ECE 411 Course Staff
//-----------------------------------------------------------------------------
// IMPORTANT: If you don't change the random seed, every time you do a `make run`
// you will run the /same/ random test. SystemVerilog calls this "random stability",
// and it's to ensure you can reproduce errors as you try to fix the DUT. Make sure
// to change the random seed or run more instructions if you want more extensive
// coverage.
//------------------------------------------------------------------------------
module random_tb
import rv32i_types::*;
(
    mem_itf_w_mask.mem itf
);

    `include "../../hvl/vcs/cp2_randinst.svh"

    RandInst gen = new();

    logic [2:0] counter;

    always_comb begin
        itf.resp[0] = 1'b1;
        itf.resp[1] = 1'b1;
    end

    // Do a bunch of LUIs to get useful register state.
    task init_register_state();
        for (int i = 0; i < 32; ++i) begin
            // @(posedge itf.clk iff |itf.rmask[0]);
            gen.randomize() with {
                instr.j_type.opcode == op_b_lui;
                instr.j_type.rd == i[4:0];
            };

            // Your code here: package these memory interactions into a task.
            itf.rdata[0] <= gen.instr.word;

            // add nops to avoid hazard
            @(posedge itf.clk iff (|itf.rmask[0]));
            itf.rdata[0] <= 32'h13;
            @(posedge itf.clk iff (|itf.rmask[0]));
            itf.rdata[0] <= 32'h13;
            @(posedge itf.clk iff (|itf.rmask[0]));
            itf.rdata[0] <= 32'h13;
            @(posedge itf.clk iff (|itf.rmask[0]));
            itf.rdata[0] <= 32'h13;
            @(posedge itf.clk iff (|itf.rmask[0]));
            itf.rdata[0] <= 32'h13;
        end
    endtask : init_register_state

    // Note that this memory model is not consistent! It ignores
    // writes and always reads out a random, valid instruction.
    task run_random_instrs();
        repeat (5000) begin
            // Always read out a valid instruction.
            if (|itf.rmask[0] || |itf.rmask[1]) begin
                if(counter == '0) begin 
                    gen.randomize() with {
                        if(instr.s_type.opcode == op_b_store) {
                            if(instr.s_type.funct3 == store_f3_sw){
                                (dut.regfile.data[instr.s_type.rs1] + instr.s_type.imm_s_bot) % 4 == 0;
                            }
                            if(instr.s_type.funct3 == store_f3_sh){
                                (dut.regfile.data[instr.s_type.rs1] + instr.s_type.imm_s_bot) % 2 == 0;
                            }
                        }
                        if(instr.i_type.opcode == op_b_load) {
                            if(instr.i_type.funct3 == load_f3_lw){
                                (dut.regfile.data[instr.i_type.rs1] + instr.i_type.i_imm) % 4 == 0;
                            }
                            if(instr.i_type.funct3 inside {load_f3_lh, load_f3_lhu}){
                                (dut.regfile.data[instr.i_type.rs1] + instr.i_type.i_imm) % 2 == 0;
                            }
                        }
                    };
                    itf.rdata[0] <= gen.instr.word;
                end else begin
                    itf.rdata[0] <= 32'h13;
                end
                counter = counter + 3'd1;
                if( counter == 3'd6 )begin
                    counter = '0;
                end
            end
        end
    endtask : run_random_instrs

    always @(posedge itf.clk iff !itf.rst) begin
        if ($isunknown(itf.rmask[0]) || $isunknown(itf.wmask[0])) begin
            $error("Memory Error: mask containes 1'bx");
            itf.error <= 1'b1;
        end
        if ((|itf.rmask[0]) && (|itf.wmask[0])) begin
            $error("Memory Error: Simultaneous memory read and write");
            itf.error <= 1'b1;
        end
        if ((|itf.rmask[0]) || (|itf.wmask[0])) begin
            if ($isunknown(itf.addr[0])) begin
                $error("Memory Error: Address contained 'x");
                itf.error <= 1'b1;
            end
            // Only check for 16-bit alignment since instructions are
            // allowed to be at 16-bit boundaries due to JALR.
            if (itf.addr[0][0] != 1'b0) begin
                $error("Memory Error: Address is not 16-bit aligned");
                itf.error <= 1'b1;
            end
        end
    end

    // A single initial block ensures random stability.
    initial begin

        // Wait for reset.
        wait(itf.rst == 1'b1);
        @(posedge itf.clk);   
        wait(itf.rst == 1'b0);

        // Get some useful state into the processor by loading in a bunch of state.
        init_register_state();
        counter = '0;
        // Run!
        run_random_instrs();

        // Finish up
        $display("Random testbench finished!");
        $finish;
    end

endmodule : random_tb
