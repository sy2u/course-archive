/home/siyingy3/Documents/ece425/mp3/pnr_workdir/pnr/regfile.lef